module cla128(a,b,ci,s,co); //single 128 bit carry lookahead adder = 32 cla4 modules
	input[127:0] a,b;
	input ci;
	output[127:0] s;
	output co;
	
	wire c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c20, c21, c22, c23, c24, c25, c26, c27, c28, c29, c30, c31;
	
	cla4 cla4_1(a[3:0],b[3:0],ci,s[3:0],c1);
	cla4 cla4_2(a[7:4],b[7:4],c1,s[7:4],c2);
	cla4 cla4_3(a[11:8],b[11:8],c2,s[11:8],c3);
	cla4 cla4_4(a[15:12],b[15:12],c3,s[15:12],c4);
	cla4 cla4_5(a[19:16],b[19:16],c4,s[19:16],c5);
	cla4 cla4_6(a[23:20],b[23:20],c5,s[23:20],c6);
	cla4 cla4_7(a[27:24],b[27:24],c6,s[27:24],c7);
	cla4 cla4_8(a[31:28],b[31:28],c7,s[31:28],c8);
	cla4 cla4_9(a[35:32],b[35:32],c8,s[35:32],c9);
	cla4 cla4_10(a[39:36],b[39:36],c9,s[39:36],c10);
	
	cla4 cla4_11(a[43:40],b[43:40],c10,s[43:40],c11);
	cla4 cla4_12(a[47:44],b[47:44],c11,s[47:44],c12);
	cla4 cla4_13(a[51:48],b[51:48],c12,s[51:48],c13);
	cla4 cla4_14(a[55:52],b[55:52],c13,s[55:52],c14);
	cla4 cla4_15(a[59:56],b[59:56],c14,s[59:56],c15);
	cla4 cla4_16(a[63:60],b[63:60],c15,s[63:60],c16);
	cla4 cla4_17(a[67:64],b[67:64],c16,s[67:64],c17);
	cla4 cla4_18(a[71:68],b[71:68],c17,s[71:68],c18);
	cla4 cla4_19(a[75:72],b[75:72],c18,s[75:72],c19);
	cla4 cla4_20(a[79:76],b[79:76],c19,s[79:76],c20);
	
	cla4 cla4_21(a[83:80],b[83:80],c20,s[83:80],c21);
	cla4 cla4_22(a[87:84],b[87:84],c21,s[87:84],c22);
	cla4 cla4_23(a[91:88],b[91:88],c22,s[91:88],c23);
	cla4 cla4_24(a[95:92],b[95:92],c23,s[95:92],c24);
	cla4 cla4_25(a[99:96],b[99:96],c24,s[99:96],c25);
	cla4 cla4_26(a[103:100],b[103:100],c25,s[103:100],c26);
	cla4 cla4_27(a[107:104],b[107:104],c26,s[107:104],c27);
	cla4 cla4_28(a[111:108],b[111:108],c27,s[111:108],c28);
	cla4 cla4_29(a[115:112],b[115:112],c28,s[115:112],c29);
	cla4 cla4_30(a[119:116],b[119:116],c29,s[119:116],c30);
	
	cla4 cla4_31(a[123:120],b[123:120],c30,s[123:120],c31);
	cla4 cla4_32(a[127:124],b[127:124],c31,s[127:124],co);
endmodule 