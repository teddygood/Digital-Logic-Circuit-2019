module _4_to_16_decoder(d, q); // 4 to 8 decoder
	input [3:0]	d; 	// select signal
	output reg [15:0] q;  
		
	always@(d)
	begin
		case(d) 
			4'b0000 : q = 16'b0000_0000_0000_0001;
			4'b0001 : q = 16'b0000_0000_0000_0010;
			4'b0010 : q = 16'b0000_0000_0000_0100;
			4'b0011 : q = 16'b0000_0000_0000_1000;
			4'b0100 : q = 16'b0000_0000_0001_0000;
			4'b0101 : q = 16'b0000_0000_0010_0000;
			4'b0110 : q = 16'b0000_0000_0100_0000;
			4'b0111 : q = 16'b0000_0000_1000_0000;
			4'b1000 : q = 16'b0000_0001_0000_0000;
			4'b1001 : q = 16'b0000_0010_0000_0000;
			4'b1010 : q = 16'b0000_0100_0000_0000;
			4'b1011 : q = 16'b0000_1000_0000_0000;
			4'b1100 : q = 16'b0001_0000_0000_0000;
			4'b1101 : q = 16'b0010_0000_0000_0000;
			4'b1110 : q = 16'b0100_0000_0000_0000;
			4'b1111 : q = 16'b1000_0000_0000_0000;
			default : q = 16'bx;
		endcase
	end
endmodule